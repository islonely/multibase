module multibase

